Daar375   17        123       Daar376   6         123       Daar377   9         123       