Daar375   17        Daar377   9         Daar376   6         